* Qucs 25.1.0  C:/Users/jnucc/Desktop/test.sch
.tran 0 10m 0.001m
.print tran v(vout)
.SUBCKT OpAmps_uA741  gnd  _net3 _net22 _net0 _net11 _net14
QT1 _net1 _net0 _net2 _net1 QMOD_T1 
.MODEL QMOD_T1 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT3 _net1 _net3 _net4 _net1 QMOD_T3 
.MODEL QMOD_T3 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT4 _net6 _net5 _net4 _net6 QMOD_T4 
.MODEL QMOD_T4 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
QT5 _net8 _net7 _net9 _net8 QMOD_T5 
.MODEL QMOD_T5 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT6 _net6 _net7 _net10 _net6 QMOD_T6 
.MODEL QMOD_T6 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT8 _net1 _net1 _net11 _net1 QMOD_T8 
.MODEL QMOD_T8 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
QT7 _net11 _net8 _net7 _net11 QMOD_T7 
.MODEL QMOD_T7 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT2 _net8 _net5 _net2 _net8 QMOD_T2 
.MODEL QMOD_T2 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
QT10 _net5 _net12 _net13 _net5 QMOD_T10 
.MODEL QMOD_T10 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT11 _net12 _net12 _net14 _net12 QMOD_T11 
.MODEL QMOD_T11 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT12 _net15 _net15 _net11 _net15 QMOD_T12 
.MODEL QMOD_T12 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
RR3 _net14 _net10 1K
RR4 _net14 _net13 5K
RR5 _net12 _net15 39K
QT9 _net5 _net1 _net11 _net5 QMOD_T9 
.MODEL QMOD_T9 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
QT14 _net16 _net6 _net17 _net16 QMOD_T14 
.MODEL QMOD_T14 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT16 _net19 _net18 _net16 _net19 QMOD_T16 
.MODEL QMOD_T16 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT17 _net16 _net17 _net20 _net16 QMOD_T17 
.MODEL QMOD_T17 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
RR6 _net19 _net18 4.5K
QT13 _net6 _net20 _net14 _net6 QMOD_T13 
.MODEL QMOD_T13 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
RR8 _net17 _net14 50K
RR9 _net20 _net14 50
RR7 _net16 _net18 7.5K
QT18 _net19 _net21 _net22 _net19 QMOD_T18 
.MODEL QMOD_T18 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT19 _net11 _net19 _net21 _net11 QMOD_T19 
.MODEL QMOD_T19 NPN(Is=2p Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
QT15 _net19 _net15 _net11 _net19 QMOD_T15 
.MODEL QMOD_T15 PNP(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=20 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
QT21 _net22 _net22 _net18 _net22 QMOD_T21 
.MODEL QMOD_T21 NPN(Is=1e-16 Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=100 Cje=3p Vje=0.75 Mje=0.33 Cjc=2p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=2p Vjs=0.75 Mjs=0 Fc=0.5 Tf=0.3n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=6n Kf=0.0 Af=1.0 Ptf=0.0) 
RR10 _net21 _net22 25
RR11 _net22 _net23 50
QT20 _net14 _net16 _net23 _net14 QMOD_T20 
.MODEL QMOD_T20 PNP(Is=2p Nf=1 Nr=1 Ikf=0 Ikr=0 Vaf=100 Var=0 Ise=0 Ne=1.5 Isc=0 Nc=2 Bf=160 Br=1 Rbm=0 Irb=0 Rc=0 Re=0 Rb=20 Cje=6p Vje=0.75 Mje=0.33 Cjc=4p Vjc=0.75 Mjc=0.33 Xcjc=1.0 Cjs=0 Vjs=0.75 Mjs=0 Fc=0.5 Tf=1n Xtf=0.0 Vtf=0.0 Itf=0.0 Tr=20n Kf=0.0 Af=1.0 Ptf=0.0) 
RR2 _net14 _net7 50K
RR1 _net14 _net9 1K
CC1 _net6 _net19 30
.ENDS

XOP1 0  _net0 _net1 volt33 volt5 0 OpAmps_uA741
XOP3 0  _net2 vout _net3 volt5 0 OpAmps_uA741
XOP2 0  _net4 _net5 volt28 volt5 0 OpAmps_uA741
R1_2 _net4 _net5  10K tc1=0.0 tc2=0.0 
R2_1 _net1 _net3  10K tc1=0.0 tc2=0.0 
R2_2 _net5 _net2  10K tc1=0.0 tc2=0.0 
R1_1 _net0 _net1  10K tc1=0.0 tc2=0.0 
R3_1 0 _net3  10K tc1=0.0 tc2=0.0 
V1 volt33 0 DC 3.3
V3 volt28 0 DC 2.8
V2 volt5 0 DC 5
RGAIN _net4 _net0  22K tc1=0.0 tc2=0.0 
R3_2 _net2 vout  10K tc1=0.0 tc2=0.0 


.END